// ----------------------------------------------------------------------
//
// File: encoder.sv
//
// Last edited: 24.07.2020
//
// Copyright (C) 2020, ETH Zurich and University of Bologna.
//
// Author: Moritz Scherer, ETH Zurich
//
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may not use this file except in compliance with the License, or, at your option, the Apache License version 2.0.
//
// You may obtain a copy of the License at
// https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//
// See the License for the specific language governing permissions and limitations under the License.
//
// ----------------------------------------------------------------------
// The encoder module is purely combinatorial and translates a 5 Trits
// to an 8-Bit tuple that is used for storage/transmission. Encoding is done in order to save storage space.
// Encodings are NOT unique, so take care.

module ternary_encoder (
                input logic [9:0]  encoder_i,
                output logic [7:0] encoder_o
                );

   logic [7:0]                     b;
   logic [9:0]                     t;

   assign encoder_o = b;
   assign t = encoder_i;

   always_comb begin

      // Optimized with Espresso for each output

      b[7] = ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[7] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & ~t[1] | t[9] & t[8] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & t[1] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | ~t[9] & ~t[8] & t[7] & t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[7] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] | t[9] & t[8] & ~t[7] & ~t[6] & ~t[5] & t[2] & t[1] & t[0] | t[9] & t[8] & t[6] & ~t[5] & t[3] & t[2] & ~t[1] & ~t[0] | t[9] & t[8] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & t[0] | ~t[9] & ~t[8] & t[7] & t[6] & ~t[5] & t[3] & t[2] & t[0] | ~t[9] & ~t[8] & t[7] & t[6] & t[5] & t[4] & t[2] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & t[3] & t[2] & ~t[1] | t[9] & t[8] & ~t[7] & t[4] & ~t[3] & ~t[2] & ~t[1] | t[9] & t[8] & ~t[7] & ~t[5] & ~t[4] & t[2] & ~t[1] | ~t[9] & ~t[8] & t[7] & t[6] & ~t[5] & ~t[3] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & ~t[3] & ~t[1] | t[9] & t[8] & t[7] & t[6] & t[4] & t[2] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & t[2] & t[0] | t[9] & t[8] & ~t[7] & ~t[5] & ~t[3] & t[0] | t[9] & t[8] & t[6] & ~t[5] & ~t[3] & ~t[1] | t[9] & t[8] & t[6] & ~t[5] & ~t[3] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[9] & t[8] & ~t[7] & t[4] & t[2] & t[0];
      b[6] = ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | t[9] & t[8] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & t[1] & t[0] | ~t[9] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | t[8] & ~t[7] & ~t[6] & t[5] & t[4] & t[3] & t[2] & t[1] & t[0] | t[8] & t[7] & t[6] & ~t[5] & ~t[3] & ~t[2] & t[1] & t[0] | ~t[9] & ~t[7] & ~t[6] & t[5] & t[4] & t[2] & t[1] & t[0] | ~t[9] & t[7] & t[6] & t[5] & t[4] & t[3] & t[2] & t[0] | t[8] & ~t[7] & ~t[6] & t[5] & t[4] & t[3] & t[2] & ~t[1] | ~t[9] & ~t[8] & t[7] & t[6] & t[5] & t[4] & t[2] & t[0] | t[8] & t[7] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & t[0] | t[8] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & ~t[1] | ~t[9] & t[7] & t[6] & t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & t[5] & t[4] & t[2] & t[0] | ~t[9] & t[7] & t[6] & t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[9] & t[8] & t[7] & t[6] & t[4] & t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & t[0] | t[8] & t[7] & t[6] & ~t[5] & ~t[3] & ~t[1] | t[8] & t[7] & t[6] & t[4] & ~t[3] & ~t[1] | t[8] & t[7] & t[6] & t[4] & ~t[3] & t[0] | t[8] & t[7] & t[6] & ~t[5] & t[2] & t[0] | t[8] & t[7] & t[6] & t[4] & t[2] & ~t[1] ;
      b[5] = ~t[9] & ~t[8] & t[7] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & ~t[1] | ~t[9] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | t[8] & ~t[7] & ~t[6] & t[5] & t[4] & t[3] & t[2] & t[1] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & ~t[7] & t[5] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[7] & ~t[6] & ~t[5] & t[3] & t[2] & t[1] & t[0] | ~t[9] & t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | ~t[9] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & t[1] & t[0] | ~t[9] & t[7] & t[6] & t[5] & t[4] & t[3] & t[2] & t[0] | t[9] & t[8] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & t[0] | ~t[9] & ~t[8] & t[7] & t[6] & ~t[5] & t[3] & t[2] & t[0] | t[8] & ~t[7] & ~t[6] & t[5] & t[4] & t[3] & t[2] & ~t[1] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] | t[9] & t[8] & t[6] & t[5] & t[4] & t[3] & t[2] & ~t[1] | ~t[9] & ~t[7] & t[5] & t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[7] & ~t[5] & ~t[4] & t[3] & t[2] & ~t[1] | t[8] & ~t[7] & ~t[6] & ~t[5] & t[3] & t[2] & ~t[1] | t[8] & ~t[7] & ~t[6] & ~t[5] & t[3] & t[2] & t[0] | ~t[9] & t[6] & t[5] & t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & t[4] & t[3] & t[2] & t[0] | ~t[9] & t[6] & t[5] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & ~t[1] | t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & ~t[3] & ~t[1] | t[8] & t[6] & t[5] & t[4] & t[2] & t[0];
      b[4] = t[9] & t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | t[9] & t[8] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & t[1] & t[0] | ~t[9] & ~t[7] & ~t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | t[8] & ~t[7] & ~t[6] & t[5] & t[4] & t[3] & t[2] & t[1] & t[0] | ~t[9] & ~t[8] & ~t[7] & t[4] & t[3] & t[2] & ~t[1] & ~t[0] | t[9] & t[8] & ~t[7] & ~t[6] & t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[7] & ~t[6] & ~t[5] & t[3] & t[2] & t[1] & t[0] | t[9] & t[8] & ~t[7] & ~t[6] & ~t[5] & t[2] & t[1] & t[0] | t[8] & t[7] & t[6] & ~t[5] & ~t[3] & ~t[2] & t[1] & t[0] | t[9] & t[8] & t[6] & ~t[5] & t[3] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[7] & ~t[6] & t[5] & t[4] & t[2] & t[1] & t[0] | ~t[9] & t[6] & t[5] & t[4] & ~t[3] & ~t[2] & t[1] & t[0] | ~t[9] & t[6] & ~t[5] & ~t[4] & t[3] & t[2] & t[1] & t[0] | t[8] & t[7] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[7] & ~t[6] & ~t[5] & ~t[3] & t[1] & t[0] | t[9] & t[8] & t[6] & t[5] & t[4] & t[3] & t[2] & ~t[1] | t[8] & ~t[7] & ~t[5] & ~t[3] & ~t[2] & t[1] & t[0] | ~t[9] & t[6] & t[4] & t[3] & t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[3] & t[1] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | t[8] & t[6] & ~t[5] & ~t[4] & t[2] & t[1] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & t[2] & t[1] & t[0] | t[8] & t[6] & t[4] & t[3] & t[2] & t[0];
      b[3] = ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[3] & t[1] & t[0] | t[8] & ~t[7] & ~t[6] & t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & t[2] & t[1] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & t[2] & ~t[1] | t[8] & t[6] & t[4] & t[2] & t[1] & t[0];
      b[2] = ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & t[0] | t[8] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[8] & t[6] & ~t[5] & ~t[4] & t[2] & t[1] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & t[0] | t[8] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] | t[8] & t[6] & t[4] & t[3] & t[2] & t[0] | t[8] & t[6] & t[4] & ~t[3] & t[0];
      b[1] = t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & t[7] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | t[8] & t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | t[8] & ~t[7] & ~t[6] & t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & t[2] & t[0] | t[8] & t[6] & ~t[5] & ~t[3] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & t[6] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & t[6] & t[4] & t[2] & t[1] & t[0] | t[8] & t[6] & t[4] & t[2] & ~t[1] ;
      b[0] = ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] & ~t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] | t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & ~t[3] & ~t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & ~t[1] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & ~t[5] & ~t[4] & t[2] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & ~t[1] | t[8] & ~t[7] & ~t[5] & ~t[3] & ~t[2] & t[1] & t[0] | ~t[9] & ~t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[8] & ~t[7] & ~t[6] & t[4] & ~t[3] & ~t[2] & t[0] | t[8] & t[6] & ~t[5] & ~t[3] & ~t[2] & t[0] | ~t[9] & ~t[8] & t[6] & t[4] & ~t[3] & ~t[2] & t[0] | ~t[9] & t[6] & t[4] & t[2] & ~t[1] & ~t[0] | t[8] & t[6] & t[4] & t[3] & t[2] & t[0] | t[8] & t[6] & t[4] & ~t[3] & t[0] | t[8] & t[6] & t[4] & t[2] & ~t[1] ;

   end // always_comb

endmodule


